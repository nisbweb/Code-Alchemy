-- Design a 2-to-1 multiplexer using VHDL. 
-- The multiplexer should take two 1-bit inputs (A and B) and a 1-bit select input (Sel).
-- The output (Y) should be A when Sel is 0, and B when Sel is 1.

-- WRITE YOUR CODE HERE