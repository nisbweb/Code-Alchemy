-- 4-bit Up/Down Counter
-- Design a 4-bit up/down counter in VHDL. 
-- The counter should count up or down based on a control signal (Up_Down), and the counting should be synchronous with the clock (Clk). 
-- The counter should reset when a reset signal (Rst) is active.

-- WRITE YOUR CODE HERE