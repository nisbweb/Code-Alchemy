-- D Flip-Flop with Asynchronous Reset
-- Design a D flip-flop with an asynchronous reset in VHDL.
-- The flip-flop should store the input D on the rising edge of the clock (Clk). If the reset (Rst) is active, the output Q should be cleared to 0, regardless of the clock.

-- WRITE YOUR CODE HERE