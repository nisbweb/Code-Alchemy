-- Parity Bit Generator
-- Design a parity bit generator in VHDL. 
-- The circuit should take an 8-bit input (Data) and output a parity bit (P) that is 1 if the number of 1s in Data is odd, and 0 if the number of 1s is even (odd parity).

-- Inputs:
-- Data: 8-bit binary input.

-- Output:
-- P: 1-bit parity output (1 for odd parity, 0 for even parity).


-- WRITE YOUR CODE HERE