-- 7-Segment Display Decoder
-- Design a 4-bit binary to 7-segment display decoder in VHDL. 
-- The decoder should take a 4-bit binary input (A) and generate the corresponding 7-segment display outputs (Seg) to display hexadecimal digits (0-9 and A-F).

-- WRITE YOUR CODE HERE
