-- Finite State Machine (FSM) for Traffic Light Controller
-- Design a finite state machine (FSM) for a traffic light controller using VHDL. 
-- The system should control a set of traffic lights with three states: Red, Yellow, and Green. The lights should transition based on a timer.

-- Inputs:
-- Clk: 1-bit clock input.
-- Rst: 1-bit reset input.

-- Outputs:
-- Red, Yellow, Green: 1-bit outputs to control the traffic lights.

-- WRITE YOUR CODE HERE